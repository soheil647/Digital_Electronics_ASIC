* Project MORB20CC
* WorkVIEW Wirelist Created with Version 3.2

X3       SRG44 N48 SHIELD44 0 BNP1S2A0
X0       5   6   N115 0 BNP2S1A1
M119     N122 0   0   0 NMOS
M120     OSGB38 OSG46 N122 0 NMOSP2
M121     VDD OSG46 OSGB38 VDD PMOSP2
X4       OSG46 N115 N38 0 BNP1S0A2
X1       N48 OS45 OS43 0 BNP1S2A0
X2       N41 OS45 N48 0 BNP1S2A0
X5       RG29 RD42 N41 0 BNP1S2A0
X6       31  N41 N38 0 BNP2S1A1


* DICTIONARY 1
* GND = 0

.GLOBAL VDD

.OPTIONS INGOLD=2 POST=2

.model NMOS
.model PMOS
.model NMOSP2
.model PMOSP2

.END
